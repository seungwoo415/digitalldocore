
.SUBCKT pass_transistors vg0 vg1 vg2 vg3 vg4 vg5 vg6 vg7 vg8 vg9 vout vdd 
 
   Xinst1 vout vg0 vdd vdd sky130_fd_pr__pfet_01v8 l=0.15u nf=1 w=0.62u
   Xinst2 vout vg1 vdd vdd sky130_fd_pr__pfet_01v8 l=0.15u nf=1 w=0.62u
   Xinst3 vout vg2 vdd vdd sky130_fd_pr__pfet_01v8 l=0.15u nf=1 w=0.62u
   Xinst4 vout vg3 vdd vdd sky130_fd_pr__pfet_01v8 l=0.15u nf=1 w=0.62u
   Xinst5 vout vg4 vdd vdd sky130_fd_pr__pfet_01v8 l=0.15u nf=1 w=0.62u
   Xinst6 vout vg5 vdd vdd sky130_fd_pr__pfet_01v8 l=0.15u nf=1 w=0.62u
   Xinst7 vout vg6 vdd vdd sky130_fd_pr__pfet_01v8 l=0.15u nf=1 w=0.62u
   Xinst8 vout vg7 vdd vdd sky130_fd_pr__pfet_01v8 l=0.15u nf=1 w=0.62u
   Xinst9 vout vg8 vdd vdd sky130_fd_pr__pfet_01v8 l=0.15u nf=1 w=0.62u
   Xinst10 vout vg9 vdd vdd sky130_fd_pr__pfet_01v8 l=0.15u nf=1 w=0.62u
 
.ENDS pass_transistors
